
`include "xcfi_macros.sv"

module xcfi_insn_spec (

    `XCFI_TRACE_INPUTS,

    `XCFI_SPEC_OUTPUTS

);

`XCFI_INSN_CHECK_COMMON

wire [63:0] insn_result = {`RS1 , `RS2} + `RS3;

assign spec_valid       = rvfi_valid && dec_xc_macc_1;
assign spec_trap        = 1'b0   ;
assign spec_rs1_addr    = `FIELD_RS1_ADDR;
assign spec_rs2_addr    = `FIELD_RS2_ADDR;
assign spec_rs3_addr    = 0;
assign spec_rd_addr     = `FIELD_RD_ADDR & 5'b11110;
assign spec_rd_wdata    = spec_rd_addr ? insn_result[31:0] : {XLEN{1'b0}};
assign spec_rd_wide     = 1'b1;
assign spec_rd_wdatahi  = insn_result[63:32];
assign spec_pc_wdata    = rvfi_pc_rdata + 4;
assign spec_mem_addr    = 0;
assign spec_mem_rmask   = 0;
assign spec_mem_wmask   = 0;
assign spec_mem_wdata   = 0;

endmodule

