`include "defines.svh"
`include "rvfi_macros.vh"

//
// module: custom_rvfi_template
//
//  A *template* module for writing custom RISC-V formal interface checkers.
//
module custom_rvfi_template (
input                                 rvfi_valid,
input  [`RISCV_FORMAL_ILEN   - 1 : 0] rvfi_insn,
input  [`RISCV_FORMAL_XLEN   - 1 : 0] rvfi_pc_rdata,
input  [`RISCV_FORMAL_XLEN   - 1 : 0] rvfi_rs1_rdata,
input  [`RISCV_FORMAL_XLEN   - 1 : 0] rvfi_rs2_rdata,
input  [`RISCV_FORMAL_XLEN   - 1 : 0] rvfi_mem_rdata,
`ifdef RISCV_FORMAL_CSR_MISA
input  [`RISCV_FORMAL_XLEN   - 1 : 0] rvfi_csr_misa_rdata,
output [`RISCV_FORMAL_XLEN   - 1 : 0] spec_csr_misa_rmask,
`endif
output                                spec_valid,
output                                spec_trap,
output [                       4 : 0] spec_rs1_addr,
output [                       4 : 0] spec_rs2_addr,
output [                       4 : 0] spec_rd_addr,
output [`RISCV_FORMAL_XLEN   - 1 : 0] spec_rd_wdata,
output [`RISCV_FORMAL_XLEN   - 1 : 0] spec_pc_wdata,
output [`RISCV_FORMAL_XLEN   - 1 : 0] spec_mem_addr,
output [`RISCV_FORMAL_XLEN/8 - 1 : 0] spec_mem_rmask,
output [`RISCV_FORMAL_XLEN/8 - 1 : 0] spec_mem_wmask,
output [`RISCV_FORMAL_XLEN   - 1 : 0] spec_mem_wdata
);

wire decoded = rvfi_valid && rvfi_insn == 32'hFFFF_FFFF;

assign spec_valid = decoded;
assign spec_trap  = 1'b1   ;

assign spec_rs1_addr = 5'd0;
assign spec_rs2_addr = 5'd0;
assign spec_rd_addr  = 5'd0;
assign spec_rd_wdata = 32'b0;
assign spec_pc_wdata = 32'b0;
assign spec_mem_rmask= 32'b0;
assign spec_mem_wmask= 32'b0;
assign spec_mem_wdata= 32'b0;

endmodule
