`define DESIGNER_ASSERTION_FETCH_BUFFER 1


